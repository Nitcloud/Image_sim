library verilog;
use verilog.vl_types.all;
entity alt_cal_mm is
    generic(
        number_of_channels: integer := 1;
        channel_address_width: integer := 1;
        sim_model_mode  : string  := "TRUE";
        lpm_type        : string  := "alt_cal_mm";
        lpm_hint        : string  := "UNUSED";
        idle            : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        ch_wait         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        testbus_set     : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi0);
        offsets_pden_rd : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        offsets_pden_wr : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi0);
        cal_pd_wr       : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi1);
        cal_rx_rd       : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi0);
        cal_rx_wr       : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi1);
        dprio_wait      : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        sample_tb       : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi1);
        test_input      : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi0);
        ch_adv          : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi0, Hi0);
        dprio_read      : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi0);
        dprio_write     : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        kick_start_rd   : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi0, Hi1);
        kick_start_wr   : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi0);
        kick_pause      : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi1);
        kick_delay_oc   : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi1, Hi0);
        sample_length   : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0)
    );
    port(
        busy            : out    vl_logic;
        cal_error       : out    vl_logic_vector;
        clock           : in     vl_logic;
        dprio_addr      : out    vl_logic_vector(15 downto 0);
        dprio_busy      : in     vl_logic;
        dprio_datain    : in     vl_logic_vector(15 downto 0);
        dprio_dataout   : out    vl_logic_vector(15 downto 0);
        dprio_rden      : out    vl_logic;
        dprio_wren      : out    vl_logic;
        quad_addr       : out    vl_logic_vector(8 downto 0);
        remap_addr      : in     vl_logic_vector(11 downto 0);
        reset           : in     vl_logic;
        retain_addr     : out    vl_logic_vector(0 downto 0);
        start           : in     vl_logic;
        transceiver_init: in     vl_logic;
        testbuses       : in     vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of number_of_channels : constant is 1;
    attribute mti_svvh_generic_type of channel_address_width : constant is 1;
    attribute mti_svvh_generic_type of sim_model_mode : constant is 1;
    attribute mti_svvh_generic_type of lpm_type : constant is 1;
    attribute mti_svvh_generic_type of lpm_hint : constant is 1;
    attribute mti_svvh_generic_type of idle : constant is 1;
    attribute mti_svvh_generic_type of ch_wait : constant is 1;
    attribute mti_svvh_generic_type of testbus_set : constant is 1;
    attribute mti_svvh_generic_type of offsets_pden_rd : constant is 1;
    attribute mti_svvh_generic_type of offsets_pden_wr : constant is 1;
    attribute mti_svvh_generic_type of cal_pd_wr : constant is 1;
    attribute mti_svvh_generic_type of cal_rx_rd : constant is 1;
    attribute mti_svvh_generic_type of cal_rx_wr : constant is 1;
    attribute mti_svvh_generic_type of dprio_wait : constant is 1;
    attribute mti_svvh_generic_type of sample_tb : constant is 1;
    attribute mti_svvh_generic_type of test_input : constant is 1;
    attribute mti_svvh_generic_type of ch_adv : constant is 1;
    attribute mti_svvh_generic_type of dprio_read : constant is 1;
    attribute mti_svvh_generic_type of dprio_write : constant is 1;
    attribute mti_svvh_generic_type of kick_start_rd : constant is 1;
    attribute mti_svvh_generic_type of kick_start_wr : constant is 1;
    attribute mti_svvh_generic_type of kick_pause : constant is 1;
    attribute mti_svvh_generic_type of kick_delay_oc : constant is 1;
    attribute mti_svvh_generic_type of sample_length : constant is 1;
end alt_cal_mm;
