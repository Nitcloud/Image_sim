library verilog;
use verilog.vl_types.all;
entity ALTERA_DEVICE_FAMILIES is
end ALTERA_DEVICE_FAMILIES;
