library verilog;
use verilog.vl_types.all;
entity altpll is
    generic(
        intended_device_family: string  := "Stratix";
        operation_mode  : string  := "NORMAL";
        pll_type        : string  := "AUTO";
        qualify_conf_done: string  := "OFF";
        compensate_clock: string  := "CLK0";
        scan_chain      : string  := "LONG";
        primary_clock   : string  := "inclk0";
        inclk0_input_frequency: integer := 1000;
        inclk1_input_frequency: integer := 0;
        gate_lock_signal: string  := "NO";
        gate_lock_counter: integer := 0;
        lock_high       : integer := 1;
        lock_low        : integer := 0;
        valid_lock_multiplier: integer := 1;
        invalid_lock_multiplier: integer := 5;
        switch_over_type: string  := "AUTO";
        switch_over_on_lossclk: string  := "OFF";
        switch_over_on_gated_lock: string  := "OFF";
        enable_switch_over_counter: string  := "OFF";
        switch_over_counter: integer := 0;
        feedback_source : string  := "EXTCLK0";
        bandwidth       : integer := 0;
        bandwidth_type  : string  := "UNUSED";
        lpm_hint        : string  := "UNUSED";
        spread_frequency: integer := 0;
        down_spread     : string  := "0.0";
        self_reset_on_gated_loss_lock: string  := "OFF";
        self_reset_on_loss_lock: string  := "OFF";
        lock_window_ui  : string  := "0.05";
        width_clock     : integer := 6;
        width_phasecounterselect: integer := 4;
        charge_pump_current_bits: integer := 9999;
        loop_filter_c_bits: integer := 9999;
        loop_filter_r_bits: integer := 9999;
        scan_chain_mif_file: string  := "UNUSED";
        simulation_type : string  := "functional";
        source_is_pll   : string  := "off";
        skip_vco        : string  := "off";
        clk9_multiply_by: integer := 1;
        clk8_multiply_by: integer := 1;
        clk7_multiply_by: integer := 1;
        clk6_multiply_by: integer := 1;
        clk5_multiply_by: integer := 1;
        clk4_multiply_by: integer := 1;
        clk3_multiply_by: integer := 1;
        clk2_multiply_by: integer := 1;
        clk1_multiply_by: integer := 1;
        clk0_multiply_by: integer := 1;
        clk9_divide_by  : integer := 1;
        clk8_divide_by  : integer := 1;
        clk7_divide_by  : integer := 1;
        clk6_divide_by  : integer := 1;
        clk5_divide_by  : integer := 1;
        clk4_divide_by  : integer := 1;
        clk3_divide_by  : integer := 1;
        clk2_divide_by  : integer := 1;
        clk1_divide_by  : integer := 1;
        clk0_divide_by  : integer := 1;
        clk9_phase_shift: string  := "0";
        clk8_phase_shift: string  := "0";
        clk7_phase_shift: string  := "0";
        clk6_phase_shift: string  := "0";
        clk5_phase_shift: string  := "0";
        clk4_phase_shift: string  := "0";
        clk3_phase_shift: string  := "0";
        clk2_phase_shift: string  := "0";
        clk1_phase_shift: string  := "0";
        clk0_phase_shift: string  := "0";
        clk5_time_delay : string  := "0";
        clk4_time_delay : string  := "0";
        clk3_time_delay : string  := "0";
        clk2_time_delay : string  := "0";
        clk1_time_delay : string  := "0";
        clk0_time_delay : string  := "0";
        clk9_duty_cycle : integer := 50;
        clk8_duty_cycle : integer := 50;
        clk7_duty_cycle : integer := 50;
        clk6_duty_cycle : integer := 50;
        clk5_duty_cycle : integer := 50;
        clk4_duty_cycle : integer := 50;
        clk3_duty_cycle : integer := 50;
        clk2_duty_cycle : integer := 50;
        clk1_duty_cycle : integer := 50;
        clk0_duty_cycle : integer := 50;
        clk9_use_even_counter_mode: string  := "OFF";
        clk8_use_even_counter_mode: string  := "OFF";
        clk7_use_even_counter_mode: string  := "OFF";
        clk6_use_even_counter_mode: string  := "OFF";
        clk5_use_even_counter_mode: string  := "OFF";
        clk4_use_even_counter_mode: string  := "OFF";
        clk3_use_even_counter_mode: string  := "OFF";
        clk2_use_even_counter_mode: string  := "OFF";
        clk1_use_even_counter_mode: string  := "OFF";
        clk0_use_even_counter_mode: string  := "OFF";
        clk9_use_even_counter_value: string  := "OFF";
        clk8_use_even_counter_value: string  := "OFF";
        clk7_use_even_counter_value: string  := "OFF";
        clk6_use_even_counter_value: string  := "OFF";
        clk5_use_even_counter_value: string  := "OFF";
        clk4_use_even_counter_value: string  := "OFF";
        clk3_use_even_counter_value: string  := "OFF";
        clk2_use_even_counter_value: string  := "OFF";
        clk1_use_even_counter_value: string  := "OFF";
        clk0_use_even_counter_value: string  := "OFF";
        clk2_output_frequency: integer := 0;
        clk1_output_frequency: integer := 0;
        clk0_output_frequency: integer := 0;
        extclk3_multiply_by: integer := 1;
        extclk2_multiply_by: integer := 1;
        extclk1_multiply_by: integer := 1;
        extclk0_multiply_by: integer := 1;
        extclk3_divide_by: integer := 1;
        extclk2_divide_by: integer := 1;
        extclk1_divide_by: integer := 1;
        extclk0_divide_by: integer := 1;
        extclk3_phase_shift: string  := "0";
        extclk2_phase_shift: string  := "0";
        extclk1_phase_shift: string  := "0";
        extclk0_phase_shift: string  := "0";
        extclk3_time_delay: string  := "0";
        extclk2_time_delay: string  := "0";
        extclk1_time_delay: string  := "0";
        extclk0_time_delay: string  := "0";
        extclk3_duty_cycle: integer := 50;
        extclk2_duty_cycle: integer := 50;
        extclk1_duty_cycle: integer := 50;
        extclk0_duty_cycle: integer := 50;
        vco_multiply_by : integer := 0;
        vco_divide_by   : integer := 0;
        sclkout0_phase_shift: string  := "0";
        sclkout1_phase_shift: string  := "0";
        dpa_multiply_by : integer := 0;
        dpa_divide_by   : integer := 0;
        dpa_divider     : integer := 0;
        vco_min         : integer := 0;
        vco_max         : integer := 0;
        vco_center      : integer := 0;
        pfd_min         : integer := 0;
        pfd_max         : integer := 0;
        m_initial       : integer := 1;
        m               : integer := 0;
        n               : integer := 1;
        m2              : integer := 1;
        n2              : integer := 1;
        ss              : integer := 0;
        l0_high         : integer := 1;
        l1_high         : integer := 1;
        g0_high         : integer := 1;
        g1_high         : integer := 1;
        g2_high         : integer := 1;
        g3_high         : integer := 1;
        e0_high         : integer := 1;
        e1_high         : integer := 1;
        e2_high         : integer := 1;
        e3_high         : integer := 1;
        l0_low          : integer := 1;
        l1_low          : integer := 1;
        g0_low          : integer := 1;
        g1_low          : integer := 1;
        g2_low          : integer := 1;
        g3_low          : integer := 1;
        e0_low          : integer := 1;
        e1_low          : integer := 1;
        e2_low          : integer := 1;
        e3_low          : integer := 1;
        l0_initial      : integer := 1;
        l1_initial      : integer := 1;
        g0_initial      : integer := 1;
        g1_initial      : integer := 1;
        g2_initial      : integer := 1;
        g3_initial      : integer := 1;
        e0_initial      : integer := 1;
        e1_initial      : integer := 1;
        e2_initial      : integer := 1;
        e3_initial      : integer := 1;
        l0_mode         : string  := "bypass";
        l1_mode         : string  := "bypass";
        g0_mode         : string  := "bypass";
        g1_mode         : string  := "bypass";
        g2_mode         : string  := "bypass";
        g3_mode         : string  := "bypass";
        e0_mode         : string  := "bypass";
        e1_mode         : string  := "bypass";
        e2_mode         : string  := "bypass";
        e3_mode         : string  := "bypass";
        l0_ph           : integer := 0;
        l1_ph           : integer := 0;
        g0_ph           : integer := 0;
        g1_ph           : integer := 0;
        g2_ph           : integer := 0;
        g3_ph           : integer := 0;
        e0_ph           : integer := 0;
        e1_ph           : integer := 0;
        e2_ph           : integer := 0;
        e3_ph           : integer := 0;
        m_ph            : integer := 0;
        l0_time_delay   : integer := 0;
        l1_time_delay   : integer := 0;
        g0_time_delay   : integer := 0;
        g1_time_delay   : integer := 0;
        g2_time_delay   : integer := 0;
        g3_time_delay   : integer := 0;
        e0_time_delay   : integer := 0;
        e1_time_delay   : integer := 0;
        e2_time_delay   : integer := 0;
        e3_time_delay   : integer := 0;
        m_time_delay    : integer := 0;
        n_time_delay    : integer := 0;
        extclk3_counter : string  := "e3";
        extclk2_counter : string  := "e2";
        extclk1_counter : string  := "e1";
        extclk0_counter : string  := "e0";
        clk9_counter    : string  := "c9";
        clk8_counter    : string  := "c8";
        clk7_counter    : string  := "c7";
        clk6_counter    : string  := "c6";
        clk5_counter    : string  := "l1";
        clk4_counter    : string  := "l0";
        clk3_counter    : string  := "g3";
        clk2_counter    : string  := "g2";
        clk1_counter    : string  := "g1";
        clk0_counter    : string  := "g0";
        enable0_counter : string  := "l0";
        enable1_counter : string  := "l0";
        charge_pump_current: integer := 2;
        loop_filter_r   : string  := "1.0";
        loop_filter_c   : integer := 5;
        vco_post_scale  : integer := 0;
        vco_frequency_control: string  := "AUTO";
        vco_phase_shift_step: integer := 0;
        lpm_type        : string  := "altpll";
        port_clkena0    : string  := "PORT_CONNECTIVITY";
        port_clkena1    : string  := "PORT_CONNECTIVITY";
        port_clkena2    : string  := "PORT_CONNECTIVITY";
        port_clkena3    : string  := "PORT_CONNECTIVITY";
        port_clkena4    : string  := "PORT_CONNECTIVITY";
        port_clkena5    : string  := "PORT_CONNECTIVITY";
        port_extclkena0 : string  := "PORT_CONNECTIVITY";
        port_extclkena1 : string  := "PORT_CONNECTIVITY";
        port_extclkena2 : string  := "PORT_CONNECTIVITY";
        port_extclkena3 : string  := "PORT_CONNECTIVITY";
        port_extclk0    : string  := "PORT_CONNECTIVITY";
        port_extclk1    : string  := "PORT_CONNECTIVITY";
        port_extclk2    : string  := "PORT_CONNECTIVITY";
        port_extclk3    : string  := "PORT_CONNECTIVITY";
        port_clk0       : string  := "PORT_CONNECTIVITY";
        port_clk1       : string  := "PORT_CONNECTIVITY";
        port_clk2       : string  := "PORT_CONNECTIVITY";
        port_clk3       : string  := "PORT_CONNECTIVITY";
        port_clk4       : string  := "PORT_CONNECTIVITY";
        port_clk5       : string  := "PORT_CONNECTIVITY";
        port_clk6       : string  := "PORT_CONNECTIVITY";
        port_clk7       : string  := "PORT_CONNECTIVITY";
        port_clk8       : string  := "PORT_CONNECTIVITY";
        port_clk9       : string  := "PORT_CONNECTIVITY";
        port_scandata   : string  := "PORT_CONNECTIVITY";
        port_scandataout: string  := "PORT_CONNECTIVITY";
        port_scandone   : string  := "PORT_CONNECTIVITY";
        port_sclkout1   : string  := "PORT_CONNECTIVITY";
        port_sclkout0   : string  := "PORT_CONNECTIVITY";
        port_clkbad0    : string  := "PORT_CONNECTIVITY";
        port_clkbad1    : string  := "PORT_CONNECTIVITY";
        port_activeclock: string  := "PORT_CONNECTIVITY";
        port_clkloss    : string  := "PORT_CONNECTIVITY";
        port_inclk1     : string  := "PORT_CONNECTIVITY";
        port_inclk0     : string  := "PORT_CONNECTIVITY";
        port_fbin       : string  := "PORT_CONNECTIVITY";
        port_fbout      : string  := "PORT_CONNECTIVITY";
        port_pllena     : string  := "PORT_CONNECTIVITY";
        port_clkswitch  : string  := "PORT_CONNECTIVITY";
        port_areset     : string  := "PORT_CONNECTIVITY";
        port_pfdena     : string  := "PORT_CONNECTIVITY";
        port_scanclk    : string  := "PORT_CONNECTIVITY";
        port_scanaclr   : string  := "PORT_CONNECTIVITY";
        port_scanread   : string  := "PORT_CONNECTIVITY";
        port_scanwrite  : string  := "PORT_CONNECTIVITY";
        port_enable0    : string  := "PORT_CONNECTIVITY";
        port_enable1    : string  := "PORT_CONNECTIVITY";
        port_locked     : string  := "PORT_CONNECTIVITY";
        port_configupdate: string  := "PORT_CONNECTIVITY";
        port_phasecounterselect: string  := "PORT_CONNECTIVITY";
        port_phasedone  : string  := "PORT_CONNECTIVITY";
        port_phasestep  : string  := "PORT_CONNECTIVITY";
        port_phaseupdown: string  := "PORT_CONNECTIVITY";
        port_vcooverrange: string  := "PORT_CONNECTIVITY";
        port_vcounderrange: string  := "PORT_CONNECTIVITY";
        port_scanclkena : string  := "PORT_CONNECTIVITY";
        using_fbmimicbidir_port: string  := "ON";
        c0_high         : integer := 1;
        c1_high         : integer := 1;
        c2_high         : integer := 1;
        c3_high         : integer := 1;
        c4_high         : integer := 1;
        c5_high         : integer := 1;
        c6_high         : integer := 1;
        c7_high         : integer := 1;
        c8_high         : integer := 1;
        c9_high         : integer := 1;
        c0_low          : integer := 1;
        c1_low          : integer := 1;
        c2_low          : integer := 1;
        c3_low          : integer := 1;
        c4_low          : integer := 1;
        c5_low          : integer := 1;
        c6_low          : integer := 1;
        c7_low          : integer := 1;
        c8_low          : integer := 1;
        c9_low          : integer := 1;
        c0_initial      : integer := 1;
        c1_initial      : integer := 1;
        c2_initial      : integer := 1;
        c3_initial      : integer := 1;
        c4_initial      : integer := 1;
        c5_initial      : integer := 1;
        c6_initial      : integer := 1;
        c7_initial      : integer := 1;
        c8_initial      : integer := 1;
        c9_initial      : integer := 1;
        c0_mode         : string  := "bypass";
        c1_mode         : string  := "bypass";
        c2_mode         : string  := "bypass";
        c3_mode         : string  := "bypass";
        c4_mode         : string  := "bypass";
        c5_mode         : string  := "bypass";
        c6_mode         : string  := "bypass";
        c7_mode         : string  := "bypass";
        c8_mode         : string  := "bypass";
        c9_mode         : string  := "bypass";
        c0_ph           : integer := 0;
        c1_ph           : integer := 0;
        c2_ph           : integer := 0;
        c3_ph           : integer := 0;
        c4_ph           : integer := 0;
        c5_ph           : integer := 0;
        c6_ph           : integer := 0;
        c7_ph           : integer := 0;
        c8_ph           : integer := 0;
        c9_ph           : integer := 0;
        c1_use_casc_in  : string  := "off";
        c2_use_casc_in  : string  := "off";
        c3_use_casc_in  : string  := "off";
        c4_use_casc_in  : string  := "off";
        c5_use_casc_in  : string  := "off";
        c6_use_casc_in  : string  := "off";
        c7_use_casc_in  : string  := "off";
        c8_use_casc_in  : string  := "off";
        c9_use_casc_in  : string  := "off";
        m_test_source   : integer := 5;
        c0_test_source  : integer := 5;
        c1_test_source  : integer := 5;
        c2_test_source  : integer := 5;
        c3_test_source  : integer := 5;
        c4_test_source  : integer := 5;
        c5_test_source  : integer := 5;
        c6_test_source  : integer := 5;
        c7_test_source  : integer := 5;
        c8_test_source  : integer := 5;
        c9_test_source  : integer := 5;
        sim_gate_lock_device_behavior: string  := "OFF"
    );
    port(
        inclk           : in     vl_logic_vector(1 downto 0);
        fbin            : in     vl_logic;
        pllena          : in     vl_logic;
        clkswitch       : in     vl_logic;
        areset          : in     vl_logic;
        pfdena          : in     vl_logic;
        clkena          : in     vl_logic_vector(5 downto 0);
        extclkena       : in     vl_logic_vector(3 downto 0);
        scanclk         : in     vl_logic;
        scanaclr        : in     vl_logic;
        scanclkena      : in     vl_logic;
        scanread        : in     vl_logic;
        scanwrite       : in     vl_logic;
        scandata        : in     vl_logic;
        phasecounterselect: in     vl_logic_vector;
        phaseupdown     : in     vl_logic;
        phasestep       : in     vl_logic;
        configupdate    : in     vl_logic;
        fbmimicbidir    : inout  vl_logic;
        clk             : out    vl_logic_vector;
        extclk          : out    vl_logic_vector(3 downto 0);
        clkbad          : out    vl_logic_vector(1 downto 0);
        enable0         : out    vl_logic;
        enable1         : out    vl_logic;
        activeclock     : out    vl_logic;
        clkloss         : out    vl_logic;
        locked          : out    vl_logic;
        scandataout     : out    vl_logic;
        scandone        : out    vl_logic;
        sclkout0        : out    vl_logic;
        sclkout1        : out    vl_logic;
        phasedone       : out    vl_logic;
        vcooverrange    : out    vl_logic;
        vcounderrange   : out    vl_logic;
        fbout           : out    vl_logic;
        fref            : out    vl_logic;
        icdrclk         : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of intended_device_family : constant is 1;
    attribute mti_svvh_generic_type of operation_mode : constant is 1;
    attribute mti_svvh_generic_type of pll_type : constant is 1;
    attribute mti_svvh_generic_type of qualify_conf_done : constant is 1;
    attribute mti_svvh_generic_type of compensate_clock : constant is 1;
    attribute mti_svvh_generic_type of scan_chain : constant is 1;
    attribute mti_svvh_generic_type of primary_clock : constant is 1;
    attribute mti_svvh_generic_type of inclk0_input_frequency : constant is 1;
    attribute mti_svvh_generic_type of inclk1_input_frequency : constant is 1;
    attribute mti_svvh_generic_type of gate_lock_signal : constant is 1;
    attribute mti_svvh_generic_type of gate_lock_counter : constant is 1;
    attribute mti_svvh_generic_type of lock_high : constant is 1;
    attribute mti_svvh_generic_type of lock_low : constant is 1;
    attribute mti_svvh_generic_type of valid_lock_multiplier : constant is 1;
    attribute mti_svvh_generic_type of invalid_lock_multiplier : constant is 1;
    attribute mti_svvh_generic_type of switch_over_type : constant is 1;
    attribute mti_svvh_generic_type of switch_over_on_lossclk : constant is 1;
    attribute mti_svvh_generic_type of switch_over_on_gated_lock : constant is 1;
    attribute mti_svvh_generic_type of enable_switch_over_counter : constant is 1;
    attribute mti_svvh_generic_type of switch_over_counter : constant is 1;
    attribute mti_svvh_generic_type of feedback_source : constant is 1;
    attribute mti_svvh_generic_type of bandwidth : constant is 1;
    attribute mti_svvh_generic_type of bandwidth_type : constant is 1;
    attribute mti_svvh_generic_type of lpm_hint : constant is 1;
    attribute mti_svvh_generic_type of spread_frequency : constant is 1;
    attribute mti_svvh_generic_type of down_spread : constant is 1;
    attribute mti_svvh_generic_type of self_reset_on_gated_loss_lock : constant is 1;
    attribute mti_svvh_generic_type of self_reset_on_loss_lock : constant is 1;
    attribute mti_svvh_generic_type of lock_window_ui : constant is 1;
    attribute mti_svvh_generic_type of width_clock : constant is 1;
    attribute mti_svvh_generic_type of width_phasecounterselect : constant is 1;
    attribute mti_svvh_generic_type of charge_pump_current_bits : constant is 1;
    attribute mti_svvh_generic_type of loop_filter_c_bits : constant is 1;
    attribute mti_svvh_generic_type of loop_filter_r_bits : constant is 1;
    attribute mti_svvh_generic_type of scan_chain_mif_file : constant is 1;
    attribute mti_svvh_generic_type of simulation_type : constant is 1;
    attribute mti_svvh_generic_type of source_is_pll : constant is 1;
    attribute mti_svvh_generic_type of skip_vco : constant is 1;
    attribute mti_svvh_generic_type of clk9_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk8_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk7_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk6_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk5_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk4_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk3_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk2_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk1_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk0_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of clk9_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk8_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk7_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk6_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk5_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk4_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk3_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk2_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk1_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk0_divide_by : constant is 1;
    attribute mti_svvh_generic_type of clk9_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk8_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk7_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk6_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk5_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk4_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk3_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk2_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk1_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk0_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of clk5_time_delay : constant is 1;
    attribute mti_svvh_generic_type of clk4_time_delay : constant is 1;
    attribute mti_svvh_generic_type of clk3_time_delay : constant is 1;
    attribute mti_svvh_generic_type of clk2_time_delay : constant is 1;
    attribute mti_svvh_generic_type of clk1_time_delay : constant is 1;
    attribute mti_svvh_generic_type of clk0_time_delay : constant is 1;
    attribute mti_svvh_generic_type of clk9_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of clk8_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of clk7_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of clk6_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of clk5_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of clk4_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of clk3_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of clk2_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of clk1_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of clk0_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of clk9_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk8_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk7_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk6_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk5_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk4_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk3_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk2_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk1_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk0_use_even_counter_mode : constant is 1;
    attribute mti_svvh_generic_type of clk9_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of clk8_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of clk7_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of clk6_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of clk5_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of clk4_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of clk3_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of clk2_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of clk1_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of clk0_use_even_counter_value : constant is 1;
    attribute mti_svvh_generic_type of clk2_output_frequency : constant is 1;
    attribute mti_svvh_generic_type of clk1_output_frequency : constant is 1;
    attribute mti_svvh_generic_type of clk0_output_frequency : constant is 1;
    attribute mti_svvh_generic_type of extclk3_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of extclk2_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of extclk1_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of extclk0_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of extclk3_divide_by : constant is 1;
    attribute mti_svvh_generic_type of extclk2_divide_by : constant is 1;
    attribute mti_svvh_generic_type of extclk1_divide_by : constant is 1;
    attribute mti_svvh_generic_type of extclk0_divide_by : constant is 1;
    attribute mti_svvh_generic_type of extclk3_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of extclk2_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of extclk1_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of extclk0_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of extclk3_time_delay : constant is 1;
    attribute mti_svvh_generic_type of extclk2_time_delay : constant is 1;
    attribute mti_svvh_generic_type of extclk1_time_delay : constant is 1;
    attribute mti_svvh_generic_type of extclk0_time_delay : constant is 1;
    attribute mti_svvh_generic_type of extclk3_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of extclk2_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of extclk1_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of extclk0_duty_cycle : constant is 1;
    attribute mti_svvh_generic_type of vco_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of vco_divide_by : constant is 1;
    attribute mti_svvh_generic_type of sclkout0_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of sclkout1_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of dpa_multiply_by : constant is 1;
    attribute mti_svvh_generic_type of dpa_divide_by : constant is 1;
    attribute mti_svvh_generic_type of dpa_divider : constant is 1;
    attribute mti_svvh_generic_type of vco_min : constant is 1;
    attribute mti_svvh_generic_type of vco_max : constant is 1;
    attribute mti_svvh_generic_type of vco_center : constant is 1;
    attribute mti_svvh_generic_type of pfd_min : constant is 1;
    attribute mti_svvh_generic_type of pfd_max : constant is 1;
    attribute mti_svvh_generic_type of m_initial : constant is 1;
    attribute mti_svvh_generic_type of m : constant is 1;
    attribute mti_svvh_generic_type of n : constant is 1;
    attribute mti_svvh_generic_type of m2 : constant is 1;
    attribute mti_svvh_generic_type of n2 : constant is 1;
    attribute mti_svvh_generic_type of ss : constant is 1;
    attribute mti_svvh_generic_type of l0_high : constant is 1;
    attribute mti_svvh_generic_type of l1_high : constant is 1;
    attribute mti_svvh_generic_type of g0_high : constant is 1;
    attribute mti_svvh_generic_type of g1_high : constant is 1;
    attribute mti_svvh_generic_type of g2_high : constant is 1;
    attribute mti_svvh_generic_type of g3_high : constant is 1;
    attribute mti_svvh_generic_type of e0_high : constant is 1;
    attribute mti_svvh_generic_type of e1_high : constant is 1;
    attribute mti_svvh_generic_type of e2_high : constant is 1;
    attribute mti_svvh_generic_type of e3_high : constant is 1;
    attribute mti_svvh_generic_type of l0_low : constant is 1;
    attribute mti_svvh_generic_type of l1_low : constant is 1;
    attribute mti_svvh_generic_type of g0_low : constant is 1;
    attribute mti_svvh_generic_type of g1_low : constant is 1;
    attribute mti_svvh_generic_type of g2_low : constant is 1;
    attribute mti_svvh_generic_type of g3_low : constant is 1;
    attribute mti_svvh_generic_type of e0_low : constant is 1;
    attribute mti_svvh_generic_type of e1_low : constant is 1;
    attribute mti_svvh_generic_type of e2_low : constant is 1;
    attribute mti_svvh_generic_type of e3_low : constant is 1;
    attribute mti_svvh_generic_type of l0_initial : constant is 1;
    attribute mti_svvh_generic_type of l1_initial : constant is 1;
    attribute mti_svvh_generic_type of g0_initial : constant is 1;
    attribute mti_svvh_generic_type of g1_initial : constant is 1;
    attribute mti_svvh_generic_type of g2_initial : constant is 1;
    attribute mti_svvh_generic_type of g3_initial : constant is 1;
    attribute mti_svvh_generic_type of e0_initial : constant is 1;
    attribute mti_svvh_generic_type of e1_initial : constant is 1;
    attribute mti_svvh_generic_type of e2_initial : constant is 1;
    attribute mti_svvh_generic_type of e3_initial : constant is 1;
    attribute mti_svvh_generic_type of l0_mode : constant is 1;
    attribute mti_svvh_generic_type of l1_mode : constant is 1;
    attribute mti_svvh_generic_type of g0_mode : constant is 1;
    attribute mti_svvh_generic_type of g1_mode : constant is 1;
    attribute mti_svvh_generic_type of g2_mode : constant is 1;
    attribute mti_svvh_generic_type of g3_mode : constant is 1;
    attribute mti_svvh_generic_type of e0_mode : constant is 1;
    attribute mti_svvh_generic_type of e1_mode : constant is 1;
    attribute mti_svvh_generic_type of e2_mode : constant is 1;
    attribute mti_svvh_generic_type of e3_mode : constant is 1;
    attribute mti_svvh_generic_type of l0_ph : constant is 1;
    attribute mti_svvh_generic_type of l1_ph : constant is 1;
    attribute mti_svvh_generic_type of g0_ph : constant is 1;
    attribute mti_svvh_generic_type of g1_ph : constant is 1;
    attribute mti_svvh_generic_type of g2_ph : constant is 1;
    attribute mti_svvh_generic_type of g3_ph : constant is 1;
    attribute mti_svvh_generic_type of e0_ph : constant is 1;
    attribute mti_svvh_generic_type of e1_ph : constant is 1;
    attribute mti_svvh_generic_type of e2_ph : constant is 1;
    attribute mti_svvh_generic_type of e3_ph : constant is 1;
    attribute mti_svvh_generic_type of m_ph : constant is 1;
    attribute mti_svvh_generic_type of l0_time_delay : constant is 1;
    attribute mti_svvh_generic_type of l1_time_delay : constant is 1;
    attribute mti_svvh_generic_type of g0_time_delay : constant is 1;
    attribute mti_svvh_generic_type of g1_time_delay : constant is 1;
    attribute mti_svvh_generic_type of g2_time_delay : constant is 1;
    attribute mti_svvh_generic_type of g3_time_delay : constant is 1;
    attribute mti_svvh_generic_type of e0_time_delay : constant is 1;
    attribute mti_svvh_generic_type of e1_time_delay : constant is 1;
    attribute mti_svvh_generic_type of e2_time_delay : constant is 1;
    attribute mti_svvh_generic_type of e3_time_delay : constant is 1;
    attribute mti_svvh_generic_type of m_time_delay : constant is 1;
    attribute mti_svvh_generic_type of n_time_delay : constant is 1;
    attribute mti_svvh_generic_type of extclk3_counter : constant is 1;
    attribute mti_svvh_generic_type of extclk2_counter : constant is 1;
    attribute mti_svvh_generic_type of extclk1_counter : constant is 1;
    attribute mti_svvh_generic_type of extclk0_counter : constant is 1;
    attribute mti_svvh_generic_type of clk9_counter : constant is 1;
    attribute mti_svvh_generic_type of clk8_counter : constant is 1;
    attribute mti_svvh_generic_type of clk7_counter : constant is 1;
    attribute mti_svvh_generic_type of clk6_counter : constant is 1;
    attribute mti_svvh_generic_type of clk5_counter : constant is 1;
    attribute mti_svvh_generic_type of clk4_counter : constant is 1;
    attribute mti_svvh_generic_type of clk3_counter : constant is 1;
    attribute mti_svvh_generic_type of clk2_counter : constant is 1;
    attribute mti_svvh_generic_type of clk1_counter : constant is 1;
    attribute mti_svvh_generic_type of clk0_counter : constant is 1;
    attribute mti_svvh_generic_type of enable0_counter : constant is 1;
    attribute mti_svvh_generic_type of enable1_counter : constant is 1;
    attribute mti_svvh_generic_type of charge_pump_current : constant is 1;
    attribute mti_svvh_generic_type of loop_filter_r : constant is 1;
    attribute mti_svvh_generic_type of loop_filter_c : constant is 1;
    attribute mti_svvh_generic_type of vco_post_scale : constant is 1;
    attribute mti_svvh_generic_type of vco_frequency_control : constant is 1;
    attribute mti_svvh_generic_type of vco_phase_shift_step : constant is 1;
    attribute mti_svvh_generic_type of lpm_type : constant is 1;
    attribute mti_svvh_generic_type of port_clkena0 : constant is 1;
    attribute mti_svvh_generic_type of port_clkena1 : constant is 1;
    attribute mti_svvh_generic_type of port_clkena2 : constant is 1;
    attribute mti_svvh_generic_type of port_clkena3 : constant is 1;
    attribute mti_svvh_generic_type of port_clkena4 : constant is 1;
    attribute mti_svvh_generic_type of port_clkena5 : constant is 1;
    attribute mti_svvh_generic_type of port_extclkena0 : constant is 1;
    attribute mti_svvh_generic_type of port_extclkena1 : constant is 1;
    attribute mti_svvh_generic_type of port_extclkena2 : constant is 1;
    attribute mti_svvh_generic_type of port_extclkena3 : constant is 1;
    attribute mti_svvh_generic_type of port_extclk0 : constant is 1;
    attribute mti_svvh_generic_type of port_extclk1 : constant is 1;
    attribute mti_svvh_generic_type of port_extclk2 : constant is 1;
    attribute mti_svvh_generic_type of port_extclk3 : constant is 1;
    attribute mti_svvh_generic_type of port_clk0 : constant is 1;
    attribute mti_svvh_generic_type of port_clk1 : constant is 1;
    attribute mti_svvh_generic_type of port_clk2 : constant is 1;
    attribute mti_svvh_generic_type of port_clk3 : constant is 1;
    attribute mti_svvh_generic_type of port_clk4 : constant is 1;
    attribute mti_svvh_generic_type of port_clk5 : constant is 1;
    attribute mti_svvh_generic_type of port_clk6 : constant is 1;
    attribute mti_svvh_generic_type of port_clk7 : constant is 1;
    attribute mti_svvh_generic_type of port_clk8 : constant is 1;
    attribute mti_svvh_generic_type of port_clk9 : constant is 1;
    attribute mti_svvh_generic_type of port_scandata : constant is 1;
    attribute mti_svvh_generic_type of port_scandataout : constant is 1;
    attribute mti_svvh_generic_type of port_scandone : constant is 1;
    attribute mti_svvh_generic_type of port_sclkout1 : constant is 1;
    attribute mti_svvh_generic_type of port_sclkout0 : constant is 1;
    attribute mti_svvh_generic_type of port_clkbad0 : constant is 1;
    attribute mti_svvh_generic_type of port_clkbad1 : constant is 1;
    attribute mti_svvh_generic_type of port_activeclock : constant is 1;
    attribute mti_svvh_generic_type of port_clkloss : constant is 1;
    attribute mti_svvh_generic_type of port_inclk1 : constant is 1;
    attribute mti_svvh_generic_type of port_inclk0 : constant is 1;
    attribute mti_svvh_generic_type of port_fbin : constant is 1;
    attribute mti_svvh_generic_type of port_fbout : constant is 1;
    attribute mti_svvh_generic_type of port_pllena : constant is 1;
    attribute mti_svvh_generic_type of port_clkswitch : constant is 1;
    attribute mti_svvh_generic_type of port_areset : constant is 1;
    attribute mti_svvh_generic_type of port_pfdena : constant is 1;
    attribute mti_svvh_generic_type of port_scanclk : constant is 1;
    attribute mti_svvh_generic_type of port_scanaclr : constant is 1;
    attribute mti_svvh_generic_type of port_scanread : constant is 1;
    attribute mti_svvh_generic_type of port_scanwrite : constant is 1;
    attribute mti_svvh_generic_type of port_enable0 : constant is 1;
    attribute mti_svvh_generic_type of port_enable1 : constant is 1;
    attribute mti_svvh_generic_type of port_locked : constant is 1;
    attribute mti_svvh_generic_type of port_configupdate : constant is 1;
    attribute mti_svvh_generic_type of port_phasecounterselect : constant is 1;
    attribute mti_svvh_generic_type of port_phasedone : constant is 1;
    attribute mti_svvh_generic_type of port_phasestep : constant is 1;
    attribute mti_svvh_generic_type of port_phaseupdown : constant is 1;
    attribute mti_svvh_generic_type of port_vcooverrange : constant is 1;
    attribute mti_svvh_generic_type of port_vcounderrange : constant is 1;
    attribute mti_svvh_generic_type of port_scanclkena : constant is 1;
    attribute mti_svvh_generic_type of using_fbmimicbidir_port : constant is 1;
    attribute mti_svvh_generic_type of c0_high : constant is 1;
    attribute mti_svvh_generic_type of c1_high : constant is 1;
    attribute mti_svvh_generic_type of c2_high : constant is 1;
    attribute mti_svvh_generic_type of c3_high : constant is 1;
    attribute mti_svvh_generic_type of c4_high : constant is 1;
    attribute mti_svvh_generic_type of c5_high : constant is 1;
    attribute mti_svvh_generic_type of c6_high : constant is 1;
    attribute mti_svvh_generic_type of c7_high : constant is 1;
    attribute mti_svvh_generic_type of c8_high : constant is 1;
    attribute mti_svvh_generic_type of c9_high : constant is 1;
    attribute mti_svvh_generic_type of c0_low : constant is 1;
    attribute mti_svvh_generic_type of c1_low : constant is 1;
    attribute mti_svvh_generic_type of c2_low : constant is 1;
    attribute mti_svvh_generic_type of c3_low : constant is 1;
    attribute mti_svvh_generic_type of c4_low : constant is 1;
    attribute mti_svvh_generic_type of c5_low : constant is 1;
    attribute mti_svvh_generic_type of c6_low : constant is 1;
    attribute mti_svvh_generic_type of c7_low : constant is 1;
    attribute mti_svvh_generic_type of c8_low : constant is 1;
    attribute mti_svvh_generic_type of c9_low : constant is 1;
    attribute mti_svvh_generic_type of c0_initial : constant is 1;
    attribute mti_svvh_generic_type of c1_initial : constant is 1;
    attribute mti_svvh_generic_type of c2_initial : constant is 1;
    attribute mti_svvh_generic_type of c3_initial : constant is 1;
    attribute mti_svvh_generic_type of c4_initial : constant is 1;
    attribute mti_svvh_generic_type of c5_initial : constant is 1;
    attribute mti_svvh_generic_type of c6_initial : constant is 1;
    attribute mti_svvh_generic_type of c7_initial : constant is 1;
    attribute mti_svvh_generic_type of c8_initial : constant is 1;
    attribute mti_svvh_generic_type of c9_initial : constant is 1;
    attribute mti_svvh_generic_type of c0_mode : constant is 1;
    attribute mti_svvh_generic_type of c1_mode : constant is 1;
    attribute mti_svvh_generic_type of c2_mode : constant is 1;
    attribute mti_svvh_generic_type of c3_mode : constant is 1;
    attribute mti_svvh_generic_type of c4_mode : constant is 1;
    attribute mti_svvh_generic_type of c5_mode : constant is 1;
    attribute mti_svvh_generic_type of c6_mode : constant is 1;
    attribute mti_svvh_generic_type of c7_mode : constant is 1;
    attribute mti_svvh_generic_type of c8_mode : constant is 1;
    attribute mti_svvh_generic_type of c9_mode : constant is 1;
    attribute mti_svvh_generic_type of c0_ph : constant is 1;
    attribute mti_svvh_generic_type of c1_ph : constant is 1;
    attribute mti_svvh_generic_type of c2_ph : constant is 1;
    attribute mti_svvh_generic_type of c3_ph : constant is 1;
    attribute mti_svvh_generic_type of c4_ph : constant is 1;
    attribute mti_svvh_generic_type of c5_ph : constant is 1;
    attribute mti_svvh_generic_type of c6_ph : constant is 1;
    attribute mti_svvh_generic_type of c7_ph : constant is 1;
    attribute mti_svvh_generic_type of c8_ph : constant is 1;
    attribute mti_svvh_generic_type of c9_ph : constant is 1;
    attribute mti_svvh_generic_type of c1_use_casc_in : constant is 1;
    attribute mti_svvh_generic_type of c2_use_casc_in : constant is 1;
    attribute mti_svvh_generic_type of c3_use_casc_in : constant is 1;
    attribute mti_svvh_generic_type of c4_use_casc_in : constant is 1;
    attribute mti_svvh_generic_type of c5_use_casc_in : constant is 1;
    attribute mti_svvh_generic_type of c6_use_casc_in : constant is 1;
    attribute mti_svvh_generic_type of c7_use_casc_in : constant is 1;
    attribute mti_svvh_generic_type of c8_use_casc_in : constant is 1;
    attribute mti_svvh_generic_type of c9_use_casc_in : constant is 1;
    attribute mti_svvh_generic_type of m_test_source : constant is 1;
    attribute mti_svvh_generic_type of c0_test_source : constant is 1;
    attribute mti_svvh_generic_type of c1_test_source : constant is 1;
    attribute mti_svvh_generic_type of c2_test_source : constant is 1;
    attribute mti_svvh_generic_type of c3_test_source : constant is 1;
    attribute mti_svvh_generic_type of c4_test_source : constant is 1;
    attribute mti_svvh_generic_type of c5_test_source : constant is 1;
    attribute mti_svvh_generic_type of c6_test_source : constant is 1;
    attribute mti_svvh_generic_type of c7_test_source : constant is 1;
    attribute mti_svvh_generic_type of c8_test_source : constant is 1;
    attribute mti_svvh_generic_type of c9_test_source : constant is 1;
    attribute mti_svvh_generic_type of sim_gate_lock_device_behavior : constant is 1;
end altpll;
